library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity GenerateurSignaux is
	
port
(
	--Entr�es
	X7_P10, X7_P9, X7_P8, X7_P7, X7_P6, X7_P5, X7_P4, X7_P3 :out std_logic;
	X6_P10, X6_P9, X6_P8, X6_P7 :out std_logic;
	S13, S14 :in std_logic; -- pour la s�lection des signaux
	Clk1M8_P18 :in std_logic
	
	--Bus
	--Bus_X7 :out std_logic_vector (0 to 7)
	--Switch :in std_logic_vector (0 to 1)
	--signaux internes
	
	
);

end GenerateurSignaux;

architecture Signaux of GenerateurSignaux is

signal Bus_X : std_logic_vector (7 downto 0); 
signal Switch : std_logic_vector (0 to 1);
signal clk4kHz : std_logic; 
signal Y 	: integer := 0; 
signal Q 	: integer := 0;  -- code par d�faut

type tab is array(0 to 239)of std_logic_vector(0 to 7);

constant Sinus 		: tab :=(x"7F",
							x"82",
							x"85",
							x"88",
							x"8C",
							x"8F",
							x"92",
							x"96",
							x"99",
							x"9C",
							x"9F",
							x"A3",
							x"A6",
							x"A9",
							x"AC",
							x"AF",
							x"B2",
							x"B5",
							x"B8",
							x"BB",
							x"BE",
							x"C1",
							x"C4",
							x"C6",
							x"C9",
							x"CC",
							x"CE",
							x"D1",
							x"D3",
							x"D6",
							x"D8",
							x"DB",
							x"DD",
							x"DF",
							x"E1",
							x"E3",
							x"E5",
							x"E7",
							x"E9",
							x"EB",
							x"EC",
							x"EE",
							x"F0",
							x"F1",
							x"F3",
							x"F4",
							x"F5",
							x"F6",
							x"F7",
							x"F8",
							x"F9",
							x"FA",
							x"FB",
							x"FB",
							x"FC",
							x"FC",
							x"FD",
							x"FD",
							x"FD",
							x"FD",
							x"FE",
							x"FD",
							x"FD",
							x"FD",
							x"FD",
							x"FC",
							x"FC",
							x"FB",
							x"FB",
							x"FA",
							x"F9",
							x"F8",
							x"F7",
							x"F6",
							x"F5",
							x"F4",
							x"F3",
							x"F1",
							x"F0",
							x"EE",
							x"EC",
							x"EB",
							x"E9",
							x"E7",
							x"E5",
							x"E3",
							x"E1",
							x"DF",
							x"DD",
							x"DB",
							x"D8",
							x"D6",
							x"D3",
							x"D1",
							x"CE",
							x"CC",
							x"C9",
							x"C6",
							x"C4",
							x"C1",
							x"BE",
							x"BB",
							x"B8",
							x"B5",
							x"B2",
							x"AF",
							x"AC",
							x"A9",
							x"A6",
							x"A3",
							x"9F",
							x"9C",
							x"99",
							x"96",
							x"92",
							x"8F",
							x"8C",
							x"88",
							x"85",
							x"82",
							x"7F",
							x"7B",
							x"78",
							x"75",
							x"71",
							x"6E",
							x"6B",
							x"67",
							x"64",
							x"61",
							x"5E",
							x"5A",
							x"57",
							x"54",
							x"51",
							x"4E",
							x"4B",
							x"48",
							x"45",
							x"42",
							x"3F",
							x"3C",
							x"39",
							x"37",
							x"34",
							x"31",
							x"2F",
							x"2C",
							x"2A",
							x"27",
							x"25",
							x"22",
							x"20",
							x"1E",
							x"1C",
							x"1A",
							x"18",
							x"16",
							x"14",
							x"12",
							x"11",
							x"0F",
							x"0D",
							x"0C",
							x"0A",
							x"09",
							x"08",
							x"07",
							x"06",
							x"05",
							x"04",
							x"03",
							x"02",
							x"02",
							x"01",
							x"01",
							x"00",
							x"00",
							x"00",
							x"00",
							x"00",
							x"00",
							x"00",
							x"00",
							x"00",
							x"01",
							x"01",
							x"02",
							x"02",
							x"03",
							x"04",
							x"05",
							x"06",
							x"07",
							x"08",
							x"09",
							x"0A",
							x"0C",
							x"0D",
							x"0F",
							x"11",
							x"12",
							x"14",
							x"16",
							x"18",
							x"1A",
							x"1C",
							x"1E",
							x"20",
							x"22",
							x"25",
							x"27",
							x"2A",
							x"2C",
							x"2F",
							x"31",
							x"34",
							x"37",
							x"39",
							x"3C",
							x"3F",
							x"42",
							x"45",
							x"48",
							x"4B",
							x"4E",
							x"51",
							x"54",
							x"57",
							x"5A",
							x"5E",
							x"61",
							x"64",
							x"67",
							x"6B",
							x"6E",
							x"71",
							x"75",
							x"78",
							x"7B"
 );
constant Sinus3		: tab :=(x"7F",
							x"88",
							x"92",
							x"9C",
							x"A6",
							x"AF",
							x"B8",
							x"C1",
							x"C9",
							x"D1",
							x"D8",
							x"DF",
							x"E5",
							x"EB",
							x"F0",
							x"F4",
							x"F7",
							x"FA",
							x"FC",
							x"FD",
							x"FE",
							x"FD",
							x"FC",
							x"FA",
							x"F7",
							x"F4",
							x"F0",
							x"EB",
							x"E5",
							x"DF",
							x"D8",
							x"D1",
							x"C9",
							x"C1",
							x"B8",
							x"AF",
							x"A6",
							x"9C",
							x"92",
							x"88",
							x"7F",
							x"75",
							x"6B",
							x"61",
							x"57",
							X"4E",
							x"45",
							x"3C",
							x"34",
							x"2C",
							x"25",
							x"1E",
							x"18",
							x"12",
							x"0D",
							x"09",
							x"06",
							x"03",
							x"01",
							x"00",
							x"00",
							x"00",
							x"01",
							x"03",
							x"06",
							x"09",
							x"0D",
							x"12",
							x"18",
							x"1E",
							x"25",
							x"2C",
							x"34",
							x"3C",
							x"45",
							x"4E",
							x"57",
							x"61",
							x"6B",
							x"75",
							x"7F",
							x"85",
							x"8C",
							x"92",
							x"98",
							x"9F",
							x"A5",
							x"AA",
							x"B0",
							x"B5",
							x"BA",
							x"BE",
							x"C2",
							x"C6",
							x"C9",
							x"CC",
							x"CE",
							x"D0",
							x"D1",
							x"D2",
							x"D3",
							x"D2",
							x"D1",
							x"D0",
							x"CE",
							x"CC",
							x"C9",
							x"C6",
							x"C2",
							x"BE",
							x"BA",
							x"B5",
							x"B0",
							x"AA",
							x"A5",
							x"9F",
							x"98",
							x"92",
							x"8C",
							x"85",
							x"7F",
							x"78",
							x"71",
							x"6B",
							x"65",
							x"5E",
							x"58",
							x"53",
							x"4D",
							x"48",
							x"43",
							x"3F",
							x"3B",
							x"37",
							x"34",
							x"31",
							x"2F",
							x"2D",
							x"2C",
							x"2B",
							x"2B",
							x"2B",
							x"2C",
							x"2D",
							x"2F",
							x"31",
							x"34",
							x"37",
							x"3B",
							x"3F",
							x"43",
							x"48",
							x"4D",
							x"53",
							x"58",
							x"5E",
							x"65",
							x"6B",
							x"71",
							x"78",
							x"7F",
							x"82",
							x"85",
							x"88",
							x"8B",
							x"8F",
							x"92",
							x"94",
							x"97",
							x"9A",
							x"9C",
							x"9E",
							x"A0",
							x"A2",
							x"A4",
							x"A5",
							x"A6",
							x"A7",
							x"A8",
							x"A8",
							x"A9",
							x"A8",
							x"A8",
							x"A7",
							x"A6",
							x"A5",
							x"A4",
							x"A2",
							x"A0",
							x"9E",
							x"9C",
							x"9A",
							x"97",
							x"94",
							x"92",
							x"8F",
							x"8B",
							x"88",
							x"85",
							x"82",
							x"7F",
							x"7B",
							x"78",
							x"75",
							x"72",
							x"6E",
							x"6B",
							x"69",
							x"66",
							x"63",
							x"61",
							x"5F",
							x"5D",
							x"5B",
							x"59",
							x"58",
							x"57",
							x"56",
							x"55",
							x"55",
							x"55",
							x"55",
							x"55",
							x"56",
							x"57",
							x"58",
							x"59",
							x"5B",
							x"5D",
							x"5F",
							x"61",
							x"63",
							x"66",
							x"69",
							x"6B",
							x"6E",
							x"72",
							x"75",
							x"78",
							x"7B"
);
constant PGTriangle	: tab :=(x"00",
							x"02",
							x"04",
							x"06",
							x"08",
							x"0A",
							x"0C",
							x"0E",
							x"10",
							x"13",
							x"15",
							x"17",
							x"19",
							x"1B",
							x"1D",
							x"1F",
							x"21",
							x"23",
							x"26",
							x"28",
							x"2A",
							x"2C",
							x"2E",
							x"30",
							x"32",
							x"34",
							x"37",
							x"39",
							x"3B",
							x"3D",
							x"3F",
							x"41",
							x"43",
							x"45",
							x"47",
							x"4A",
							x"4C",
							x"4E",
							x"50",
							x"52",
							x"54",
							x"56",
							x"58",
							x"5B",
							x"5D",
							x"5F",
							x"61",
							x"63",
							x"65",
							x"67",
							x"69",
							x"6B",
							x"6E",
							x"70",
							x"72",
							x"74",
							x"76",
							x"78",
							x"7A",
							x"7C",
							x"7F",
							x"7C",
							x"7A",
							x"78",
							x"76",
							x"74",
							x"72",
							x"70",
							x"6E",
							x"6B",
							x"69",
							x"67",
							x"65",
							x"63",
							x"61",
							x"5F",
							x"5D",
							x"5B",
							x"58",
							x"56",
							x"54",
							x"52",
							x"50",
							x"4E",
							x"4C",
							x"4A",
							x"47",
							x"45",
							x"43",
							x"41",
							x"3F",
							x"3D",
							x"3B",
							x"39",
							x"37",
							x"34",
							x"32",
							x"30",
							x"2E",
							x"2C",
							x"2A",
							x"28",
							x"26",
							x"23",
							x"21",
							x"1F",
							x"1D",
							x"1B",
							x"19",
							x"17",
							x"15",
							x"13",
							x"10",
							x"0E",
							x"0C",
							x"0A",
							x"08",
							x"06",
							x"04",
							x"02",
							x"00",
							x"04",
							x"08",
							x"0C",
							x"11",
							x"15",
							x"19",
							x"1D",
							x"22",
							x"26",
							x"2A",
							x"2E",
							x"33",
							x"37",
							x"3B",
							x"3F",
							x"44",
							x"48",
							x"4C",
							x"50",
							x"55",
							x"59",
							x"5D",
							x"61",
							x"66",
							x"6A",
							x"6E",
							x"72",
							x"77",
							x"7B",
							x"7F",
							x"83",
							x"88",
							x"8C",
							x"90",
							x"94",
							x"99",
							x"9D",
							x"A1",
							x"A5",
							x"AA",
							x"AE",
							x"B2",
							x"B6",
							x"BB",
							x"BF",
							x"C3",
							x"C7",
							x"CC",
							x"D0",
							x"D4",
							x"D8",
							x"DD",
							x"E1",
							x"E5",
							x"E9",
							x"EE",
							x"F2",
							x"F6",
							x"FA",
							x"FF",
							x"FA",
							x"F6",
							x"F2",
							x"EE",
							x"E9",
							x"E5",
							x"E1",
							x"DD",
							x"D8",
							x"D4",
							x"D0",
							x"CC",
							x"C7",
							x"C3",
							x"BF",
							x"BB",
							x"B6",
							x"B2",
							x"AE",
							x"AA",
							x"A5",
							x"A1",
							x"9D",
							x"99",
							x"94",
							x"90",
							x"8C",
							x"88",
							x"83",
							x"7F",
							x"7B",
							x"77",
							x"72",
							x"6E",
							x"6A",
							x"66",
							x"61",
							x"5D",
							x"59",
							x"55",
							x"50",
							x"4C",
							x"48",
							x"44",
							x"3F",
							x"3B",
							x"37",
							x"33",
							x"2E",
							x"2A",
							x"26",
							x"22",
							x"1D",
							x"19",
							x"15",
							x"11",
							x"0C",
							x"08",
							x"04"
							);
constant Triangle3 	: tab :=(x"00",
							x"03",
							x"06",
							x"09",
							x"0C",
							x"0F",
							x"13",
							x"16",
							x"19",
							x"1C",
							x"1F",
							x"22",
							x"26",
							x"29",
							x"2C",
							x"2F",
							x"32",
							x"35",
							x"39",
							x"3C",
							x"3F",
							x"42",
							x"45",
							x"49",
							x"4C",
							x"4F",
							x"52",
							x"55",
							x"58",
							x"5C",
							x"5F",
							x"62",
							x"65",
							x"68",
							x"6B",
							x"6F",
							x"72",
							x"75",
							x"78",
							x"7B",
							x"7F",
							x"7B",
							x"78",
							x"75",
							x"72",
							x"6F",
							x"6B",
							x"68",
							x"65",
							x"62",
							x"5F",
							x"5C",
							x"58",
							x"55",
							x"52",
							x"4F",
							x"4C",
							x"49",
							x"45",
							x"42",
							x"3F",
							x"3C",
							x"39",
							x"35",
							x"32",
							x"2F",
							x"2C",
							x"29",
							x"26",
							x"22",
							x"1F",
							x"1C",
							x"19",
							x"16",
							x"13",
							x"0F",
							x"0C",
							x"09",
							x"06",
							x"03",
							x"00",
							x"06",
							x"0C",
							x"13",
							x"19",
							x"1F",
							x"26",
							x"2C",
							x"33",
							x"39",
							x"3F",
							x"46",
							x"4C",
							x"52",
							x"59",
							x"5F",
							x"66",
							x"6C",
							x"72",
							x"79",
							x"7F",
							x"85",
							x"8C",
							x"92",
							x"99",
							x"9F",
							x"A5",
							x"AC",
							x"B2",
							x"B8",
							x"BF",
							x"C5",
							x"CC",
							x"D2",
							x"D8",
							x"DF",
							x"E5",
							x"EB",
							x"F2",
							x"F8",
							x"FF",
							x"F8",
							x"F2",
							x"EB",
							x"E5",
							x"DF",
							x"D8",
							x"D2",
							x"CC",
							x"C5",
							x"BF",
							x"B8",
							x"B2",
							x"AC",
							x"A5",
							x"9F",
							x"99",
							x"92",
							x"8C",
							x"85",
							x"7F",
							x"79",
							x"72",
							x"6C",
							x"66",
							x"5F",
							x"59",
							x"52",
							x"4C",
							x"46",
							x"3F",
							x"39",
							x"33",
							x"2C",
							x"26",
							x"1F",
							x"19",
							x"13",
							x"0C",
							x"06",
							x"00",
							x"03",
							x"06",
							x"09",
							x"0C",
							x"0F",
							x"13",
							x"16",
							x"19",
							x"1C",
							x"1F",
							x"22",
							x"26",
							x"29",
							x"2C",
							x"2F",
							x"32",
							x"35",
							x"39",
							x"3C",
							x"3F",
							x"42",
							x"45",
							x"49",
							x"4C",
							x"4F",
							x"52",
							x"55",
							x"58",
							x"5C",
							x"5F",
							x"62",
							x"65",
							x"68",
							x"6B",
							x"6F",
							x"72",
							x"75",
							x"78",
							x"7B",
							x"7F",
							x"7B",
							x"78",
							x"75",
							x"72",
							x"6F",
							x"6B",
							x"68",
							x"65",
							x"62",
							x"5F",
							x"5C",
							x"58",
							x"55",
							x"52",
							x"4F",
							x"4C",
							x"49",
							x"45",
							x"42",
							x"3F",
							x"3C",
							x"39",
							x"35",
							x"32",
							x"2F",
							x"2C",
							x"29",
							x"26",
							x"22",
							x"1F",
							x"1C",
							x"19",
							x"16",
							x"13",
							x"0F",
							x"0C",
							x"09",
							x"06",
							x"03"
							);
begin 
	--Bus_X <= (X7_P10, X7_P9, X7_P8, X7_P7, X7_P6, X7_P5, X7_P4, X7_P3);
	X7_P10 <= Bus_X(0); 
	X7_P9 <= Bus_X(1);
	X7_P8 <= Bus_X(2);
	X7_P7 <= Bus_X(3);
	X7_P6 <= Bus_X(4);
	X7_P5 <= Bus_X(5);
	X7_P4 <= Bus_X(6);
	X7_P3 <= Bus_X(7);
	Switch<=(S13,S14);	
	

	--Switch <= (S13, S14);
	main : process(clk4kHz) 
		begin
		X6_P8	<= '0';
		X6_P9	<= '0';
		X6_P10	<= '1';
		if rising_edge (clk4kHz) then
			if Y >= 240 then
				Y <= 0;
			else
				Y <= Y+1;
			end if;
		end if;
			case Switch is
				when "00" => Bus_X <= Sinus(Y);
				when "01" => Bus_X <= Sinus3(Y);
				when "10" => Bus_X <= PGTriangle(Y);
				when "11" => Bus_X <= Triangle3(Y);
			end case;
	end process;			
		clock:process (Clk1M8_P18)
		begin
			if rising_edge(Clk1M8_P18)then
				if Q >= 920 then				--division du quartz de 1,8MHz (4kHz)
					Q <= 0;
					if clk4kHz = '0' then			
						clk4kHz <= '1';
						X6_P7	<= '0';
												
					else 
						clk4kHz <= '0';
						X6_P7	<= '1';

					end if; 					
			    else
					Q <= Q +1;	
				end if;		
			end if;
			
		end process;
end Signaux;